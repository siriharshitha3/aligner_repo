///////////////////////////////////////////////////////////////////////////////
// File:        cfs_apb_sequence_rw.sv
// Author:      Cristian Florin Slav
// Date:        2023-08-23
// Description: APB read-write sequence class.
///////////////////////////////////////////////////////////////////////////////
`ifndef CFS_APB_SEQUENCE_RW_SV
  `define CFS_APB_SEQUENCE_RW_SV

  class cfs_apb_sequence_rw extends cfs_apb_sequence_base;
    
    //Address
    rand cfs_apb_addr addr;
    
    //Write data
    rand cfs_apb_data wr_data;
    
    `uvm_object_utils(cfs_apb_sequence_rw)
    
    function new(string name = "");
      super.new(name);
    endfunction
    
    virtual task body();
//       cfs_apb_item_drv item = cfs_apb_item_drv::type_id::create("item");
      
//       void'(item.randomize() with {
//         dir  == CFS_APB_READ;
//         //Pay attention to the "local::" in order to avoid name confusion
//         addr == local::addr;
//       });
//       start_item(item);
//       finish_item(item);
      
//       void'(item.randomize() with {
//         dir  == CFS_APB_WRITE;
//         //Pay attention to the "local::" in order to avoid name confusion
//         addr == local::addr;
//         data == wr_data;
//       });
//       start_item(item);
//       finish_item(item);
      
      //The above code can be replaced with `uvm_do macros
      cfs_apb_item_drv item;
      
      `uvm_do_with(item, {
        dir  == CFS_APB_READ;
        addr == local::addr;
      });
      
      `uvm_do_with(item, {
        dir  == CFS_APB_WRITE;
        addr == local::addr;
        data == wr_data;
      });
      
    endtask

  endclass

`endif